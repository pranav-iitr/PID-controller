`timescale 1ns / 1ps
module multiplier(m1,m2,out);
input[15:0] m1; 
input[15:0] m2; 
output[15:0] out; 
wire [31:0]M;
wire m1m2_00;
wire m1m2_01;
wire m1m2_02;
wire m1m2_03;
wire m1m2_04;
wire m1m2_05;
wire m1m2_06;
wire m1m2_07;
wire m1m2_08;
wire m1m2_09;
wire m1m2_010;
wire m1m2_011;
wire m1m2_012;
wire m1m2_013;
wire m1m2_014;
wire m1m2_015;
wire m1m2_10;
wire m1m2_11;
wire m1m2_12;
wire m1m2_13;
wire m1m2_14;
wire m1m2_15;
wire m1m2_16;
wire m1m2_17;
wire m1m2_18;
wire m1m2_19;
wire m1m2_110;
wire m1m2_111;
wire m1m2_112;
wire m1m2_113;
wire m1m2_114;
wire m1m2_115;
wire m1m2_20;
wire m1m2_21;
wire m1m2_22;
wire m1m2_23;
wire m1m2_24;
wire m1m2_25;
wire m1m2_26;
wire m1m2_27;
wire m1m2_28;
wire m1m2_29;
wire m1m2_210;
wire m1m2_211;
wire m1m2_212;
wire m1m2_213;
wire m1m2_214;
wire m1m2_215;
wire m1m2_30;
wire m1m2_31;
wire m1m2_32;
wire m1m2_33;
wire m1m2_34;
wire m1m2_35;
wire m1m2_36;
wire m1m2_37;
wire m1m2_38;
wire m1m2_39;
wire m1m2_310;
wire m1m2_311;
wire m1m2_312;
wire m1m2_313;
wire m1m2_314;
wire m1m2_315;
wire m1m2_40;
wire m1m2_41;
wire m1m2_42;
wire m1m2_43;
wire m1m2_44;
wire m1m2_45;
wire m1m2_46;
wire m1m2_47;
wire m1m2_48;
wire m1m2_49;
wire m1m2_410;
wire m1m2_411;
wire m1m2_412;
wire m1m2_413;
wire m1m2_414;
wire m1m2_415;
wire m1m2_50;
wire m1m2_51;
wire m1m2_52;
wire m1m2_53;
wire m1m2_54;
wire m1m2_55;
wire m1m2_56;
wire m1m2_57;
wire m1m2_58;
wire m1m2_59;
wire m1m2_510;
wire m1m2_511;
wire m1m2_512;
wire m1m2_513;
wire m1m2_514;
wire m1m2_515;
wire m1m2_60;
wire m1m2_61;
wire m1m2_62;
wire m1m2_63;
wire m1m2_64;
wire m1m2_65;
wire m1m2_66;
wire m1m2_67;
wire m1m2_68;
wire m1m2_69;
wire m1m2_610;
wire m1m2_611;
wire m1m2_612;
wire m1m2_613;
wire m1m2_614;
wire m1m2_615;
wire m1m2_70;
wire m1m2_71;
wire m1m2_72;
wire m1m2_73;
wire m1m2_74;
wire m1m2_75;
wire m1m2_76;
wire m1m2_77;
wire m1m2_78;
wire m1m2_79;
wire m1m2_710;
wire m1m2_711;
wire m1m2_712;
wire m1m2_713;
wire m1m2_714;
wire m1m2_715;
wire m1m2_80;
wire m1m2_81;
wire m1m2_82;
wire m1m2_83;
wire m1m2_84;
wire m1m2_85;
wire m1m2_86;
wire m1m2_87;
wire m1m2_88;
wire m1m2_89;
wire m1m2_810;
wire m1m2_811;
wire m1m2_812;
wire m1m2_813;
wire m1m2_814;
wire m1m2_815;
wire m1m2_90;
wire m1m2_91;
wire m1m2_92;
wire m1m2_93;
wire m1m2_94;
wire m1m2_95;
wire m1m2_96;
wire m1m2_97;
wire m1m2_98;
wire m1m2_99;
wire m1m2_910;
wire m1m2_911;
wire m1m2_912;
wire m1m2_913;
wire m1m2_914;
wire m1m2_915;
wire m1m2_100;
wire m1m2_101;
wire m1m2_102;
wire m1m2_103;
wire m1m2_104;
wire m1m2_105;
wire m1m2_106;
wire m1m2_107;
wire m1m2_108;
wire m1m2_109;
wire m1m2_1010;
wire m1m2_1011;
wire m1m2_1012;
wire m1m2_1013;
wire m1m2_1014;
wire m1m2_1015;
wire m1m2_110;
wire m1m2_111;
wire m1m2_112;
wire m1m2_113;
wire m1m2_114;
wire m1m2_115;
wire m1m2_116;
wire m1m2_117;
wire m1m2_118;
wire m1m2_119;
wire m1m2_1110;
wire m1m2_1111;
wire m1m2_1112;
wire m1m2_1113;
wire m1m2_1114;
wire m1m2_1115;
wire m1m2_120;
wire m1m2_121;
wire m1m2_122;
wire m1m2_123;
wire m1m2_124;
wire m1m2_125;
wire m1m2_126;
wire m1m2_127;
wire m1m2_128;
wire m1m2_129;
wire m1m2_1210;
wire m1m2_1211;
wire m1m2_1212;
wire m1m2_1213;
wire m1m2_1214;
wire m1m2_1215;
wire m1m2_130;
wire m1m2_131;
wire m1m2_132;
wire m1m2_133;
wire m1m2_134;
wire m1m2_135;
wire m1m2_136;
wire m1m2_137;
wire m1m2_138;
wire m1m2_139;
wire m1m2_1310;
wire m1m2_1311;
wire m1m2_1312;
wire m1m2_1313;
wire m1m2_1314;
wire m1m2_1315;
wire m1m2_140;
wire m1m2_141;
wire m1m2_142;
wire m1m2_143;
wire m1m2_144;
wire m1m2_145;
wire m1m2_146;
wire m1m2_147;
wire m1m2_148;
wire m1m2_149;
wire m1m2_1410;
wire m1m2_1411;
wire m1m2_1412;
wire m1m2_1413;
wire m1m2_1414;
wire m1m2_1415;
wire m1m2_150;
wire m1m2_151;
wire m1m2_152;
wire m1m2_153;
wire m1m2_154;
wire m1m2_155;
wire m1m2_156;
wire m1m2_157;
wire m1m2_158;
wire m1m2_159;
wire m1m2_1510;
wire m1m2_1511;
wire m1m2_1512;
wire m1m2_1513;
wire m1m2_1514;
wire m1m2_1515;
wire[15:0] p0;
wire[15:0] sum1;
wire c1;
wire[15:0] p1;
wire[15:0] sum2;
wire c2;
wire[15:0] p2;
wire[15:0] sum3;
wire c3;
wire[15:0] p3;
wire[15:0] sum4;
wire c4;
wire[15:0] p4;
wire[15:0] sum5;
wire c5;
wire[15:0] p5;
wire[15:0] sum6;
wire c6;
wire[15:0] p6;
wire[15:0] sum7;
wire c7;
wire[15:0] p7;
wire[15:0] sum8;
wire c8;
wire[15:0] p8;
wire[15:0] sum9;
wire c9;
wire[15:0] p9;
wire[15:0] sum10;
wire c10;
wire[15:0] p10;
wire[15:0] sum11;
wire c11;
wire[15:0] p11;
wire[15:0] sum12;
wire c12;
wire[15:0] p12;
wire[15:0] sum13;
wire c13;
wire[15:0] p13;
wire[15:0] sum14;
wire c14;
wire[15:0] p14;
wire[15:0] sum15;
wire c15;
wire[15:0] p15;
and(m1m2_00,m1[0],m2[0]);
and(m1m2_01,m1[0],m2[1]);
and(m1m2_02,m1[0],m2[2]);
and(m1m2_03,m1[0],m2[3]);
and(m1m2_04,m1[0],m2[4]);
and(m1m2_05,m1[0],m2[5]);
and(m1m2_06,m1[0],m2[6]);
and(m1m2_07,m1[0],m2[7]);
and(m1m2_08,m1[0],m2[8]);
and(m1m2_09,m1[0],m2[9]);
and(m1m2_010,m1[0],m2[10]);
and(m1m2_011,m1[0],m2[11]);
and(m1m2_012,m1[0],m2[12]);
and(m1m2_013,m1[0],m2[13]);
and(m1m2_014,m1[0],m2[14]);
and(m1m2_015,m1[0],m2[15]);
and(m1m2_10,m1[1],m2[0]);
and(m1m2_11,m1[1],m2[1]);
and(m1m2_12,m1[1],m2[2]);
and(m1m2_13,m1[1],m2[3]);
and(m1m2_14,m1[1],m2[4]);
and(m1m2_15,m1[1],m2[5]);
and(m1m2_16,m1[1],m2[6]);
and(m1m2_17,m1[1],m2[7]);
and(m1m2_18,m1[1],m2[8]);
and(m1m2_19,m1[1],m2[9]);
and(m1m2_110,m1[1],m2[10]);
and(m1m2_111,m1[1],m2[11]);
and(m1m2_112,m1[1],m2[12]);
and(m1m2_113,m1[1],m2[13]);
and(m1m2_114,m1[1],m2[14]);
and(m1m2_115,m1[1],m2[15]);
and(m1m2_20,m1[2],m2[0]);
and(m1m2_21,m1[2],m2[1]);
and(m1m2_22,m1[2],m2[2]);
and(m1m2_23,m1[2],m2[3]);
and(m1m2_24,m1[2],m2[4]);
and(m1m2_25,m1[2],m2[5]);
and(m1m2_26,m1[2],m2[6]);
and(m1m2_27,m1[2],m2[7]);
and(m1m2_28,m1[2],m2[8]);
and(m1m2_29,m1[2],m2[9]);
and(m1m2_210,m1[2],m2[10]);
and(m1m2_211,m1[2],m2[11]);
and(m1m2_212,m1[2],m2[12]);
and(m1m2_213,m1[2],m2[13]);
and(m1m2_214,m1[2],m2[14]);
and(m1m2_215,m1[2],m2[15]);
and(m1m2_30,m1[3],m2[0]);
and(m1m2_31,m1[3],m2[1]);
and(m1m2_32,m1[3],m2[2]);
and(m1m2_33,m1[3],m2[3]);
and(m1m2_34,m1[3],m2[4]);
and(m1m2_35,m1[3],m2[5]);
and(m1m2_36,m1[3],m2[6]);
and(m1m2_37,m1[3],m2[7]);
and(m1m2_38,m1[3],m2[8]);
and(m1m2_39,m1[3],m2[9]);
and(m1m2_310,m1[3],m2[10]);
and(m1m2_311,m1[3],m2[11]);
and(m1m2_312,m1[3],m2[12]);
and(m1m2_313,m1[3],m2[13]);
and(m1m2_314,m1[3],m2[14]);
and(m1m2_315,m1[3],m2[15]);
and(m1m2_40,m1[4],m2[0]);
and(m1m2_41,m1[4],m2[1]);
and(m1m2_42,m1[4],m2[2]);
and(m1m2_43,m1[4],m2[3]);
and(m1m2_44,m1[4],m2[4]);
and(m1m2_45,m1[4],m2[5]);
and(m1m2_46,m1[4],m2[6]);
and(m1m2_47,m1[4],m2[7]);
and(m1m2_48,m1[4],m2[8]);
and(m1m2_49,m1[4],m2[9]);
and(m1m2_410,m1[4],m2[10]);
and(m1m2_411,m1[4],m2[11]);
and(m1m2_412,m1[4],m2[12]);
and(m1m2_413,m1[4],m2[13]);
and(m1m2_414,m1[4],m2[14]);
and(m1m2_415,m1[4],m2[15]);
and(m1m2_50,m1[5],m2[0]);
and(m1m2_51,m1[5],m2[1]);
and(m1m2_52,m1[5],m2[2]);
and(m1m2_53,m1[5],m2[3]);
and(m1m2_54,m1[5],m2[4]);
and(m1m2_55,m1[5],m2[5]);
and(m1m2_56,m1[5],m2[6]);
and(m1m2_57,m1[5],m2[7]);
and(m1m2_58,m1[5],m2[8]);
and(m1m2_59,m1[5],m2[9]);
and(m1m2_510,m1[5],m2[10]);
and(m1m2_511,m1[5],m2[11]);
and(m1m2_512,m1[5],m2[12]);
and(m1m2_513,m1[5],m2[13]);
and(m1m2_514,m1[5],m2[14]);
and(m1m2_515,m1[5],m2[15]);
and(m1m2_60,m1[6],m2[0]);
and(m1m2_61,m1[6],m2[1]);
and(m1m2_62,m1[6],m2[2]);
and(m1m2_63,m1[6],m2[3]);
and(m1m2_64,m1[6],m2[4]);
and(m1m2_65,m1[6],m2[5]);
and(m1m2_66,m1[6],m2[6]);
and(m1m2_67,m1[6],m2[7]);
and(m1m2_68,m1[6],m2[8]);
and(m1m2_69,m1[6],m2[9]);
and(m1m2_610,m1[6],m2[10]);
and(m1m2_611,m1[6],m2[11]);
and(m1m2_612,m1[6],m2[12]);
and(m1m2_613,m1[6],m2[13]);
and(m1m2_614,m1[6],m2[14]);
and(m1m2_615,m1[6],m2[15]);
and(m1m2_70,m1[7],m2[0]);
and(m1m2_71,m1[7],m2[1]);
and(m1m2_72,m1[7],m2[2]);
and(m1m2_73,m1[7],m2[3]);
and(m1m2_74,m1[7],m2[4]);
and(m1m2_75,m1[7],m2[5]);
and(m1m2_76,m1[7],m2[6]);
and(m1m2_77,m1[7],m2[7]);
and(m1m2_78,m1[7],m2[8]);
and(m1m2_79,m1[7],m2[9]);
and(m1m2_710,m1[7],m2[10]);
and(m1m2_711,m1[7],m2[11]);
and(m1m2_712,m1[7],m2[12]);
and(m1m2_713,m1[7],m2[13]);
and(m1m2_714,m1[7],m2[14]);
and(m1m2_715,m1[7],m2[15]);
and(m1m2_80,m1[8],m2[0]);
and(m1m2_81,m1[8],m2[1]);
and(m1m2_82,m1[8],m2[2]);
and(m1m2_83,m1[8],m2[3]);
and(m1m2_84,m1[8],m2[4]);
and(m1m2_85,m1[8],m2[5]);
and(m1m2_86,m1[8],m2[6]);
and(m1m2_87,m1[8],m2[7]);
and(m1m2_88,m1[8],m2[8]);
and(m1m2_89,m1[8],m2[9]);
and(m1m2_810,m1[8],m2[10]);
and(m1m2_811,m1[8],m2[11]);
and(m1m2_812,m1[8],m2[12]);
and(m1m2_813,m1[8],m2[13]);
and(m1m2_814,m1[8],m2[14]);
and(m1m2_815,m1[8],m2[15]);
and(m1m2_90,m1[9],m2[0]);
and(m1m2_91,m1[9],m2[1]);
and(m1m2_92,m1[9],m2[2]);
and(m1m2_93,m1[9],m2[3]);
and(m1m2_94,m1[9],m2[4]);
and(m1m2_95,m1[9],m2[5]);
and(m1m2_96,m1[9],m2[6]);
and(m1m2_97,m1[9],m2[7]);
and(m1m2_98,m1[9],m2[8]);
and(m1m2_99,m1[9],m2[9]);
and(m1m2_910,m1[9],m2[10]);
and(m1m2_911,m1[9],m2[11]);
and(m1m2_912,m1[9],m2[12]);
and(m1m2_913,m1[9],m2[13]);
and(m1m2_914,m1[9],m2[14]);
and(m1m2_915,m1[9],m2[15]);
and(m1m2_100,m1[10],m2[0]);
and(m1m2_101,m1[10],m2[1]);
and(m1m2_102,m1[10],m2[2]);
and(m1m2_103,m1[10],m2[3]);
and(m1m2_104,m1[10],m2[4]);
and(m1m2_105,m1[10],m2[5]);
and(m1m2_106,m1[10],m2[6]);
and(m1m2_107,m1[10],m2[7]);
and(m1m2_108,m1[10],m2[8]);
and(m1m2_109,m1[10],m2[9]);
and(m1m2_1010,m1[10],m2[10]);
and(m1m2_1011,m1[10],m2[11]);
and(m1m2_1012,m1[10],m2[12]);
and(m1m2_1013,m1[10],m2[13]);
and(m1m2_1014,m1[10],m2[14]);
and(m1m2_1015,m1[10],m2[15]);
and(m1m2_110,m1[11],m2[0]);
and(m1m2_111,m1[11],m2[1]);
and(m1m2_112,m1[11],m2[2]);
and(m1m2_113,m1[11],m2[3]);
and(m1m2_114,m1[11],m2[4]);
and(m1m2_115,m1[11],m2[5]);
and(m1m2_116,m1[11],m2[6]);
and(m1m2_117,m1[11],m2[7]);
and(m1m2_118,m1[11],m2[8]);
and(m1m2_119,m1[11],m2[9]);
and(m1m2_1110,m1[11],m2[10]);
and(m1m2_1111,m1[11],m2[11]);
and(m1m2_1112,m1[11],m2[12]);
and(m1m2_1113,m1[11],m2[13]);
and(m1m2_1114,m1[11],m2[14]);
and(m1m2_1115,m1[11],m2[15]);
and(m1m2_120,m1[12],m2[0]);
and(m1m2_121,m1[12],m2[1]);
and(m1m2_122,m1[12],m2[2]);
and(m1m2_123,m1[12],m2[3]);
and(m1m2_124,m1[12],m2[4]);
and(m1m2_125,m1[12],m2[5]);
and(m1m2_126,m1[12],m2[6]);
and(m1m2_127,m1[12],m2[7]);
and(m1m2_128,m1[12],m2[8]);
and(m1m2_129,m1[12],m2[9]);
and(m1m2_1210,m1[12],m2[10]);
and(m1m2_1211,m1[12],m2[11]);
and(m1m2_1212,m1[12],m2[12]);
and(m1m2_1213,m1[12],m2[13]);
and(m1m2_1214,m1[12],m2[14]);
and(m1m2_1215,m1[12],m2[15]);
and(m1m2_130,m1[13],m2[0]);
and(m1m2_131,m1[13],m2[1]);
and(m1m2_132,m1[13],m2[2]);
and(m1m2_133,m1[13],m2[3]);
and(m1m2_134,m1[13],m2[4]);
and(m1m2_135,m1[13],m2[5]);
and(m1m2_136,m1[13],m2[6]);
and(m1m2_137,m1[13],m2[7]);
and(m1m2_138,m1[13],m2[8]);
and(m1m2_139,m1[13],m2[9]);
and(m1m2_1310,m1[13],m2[10]);
and(m1m2_1311,m1[13],m2[11]);
and(m1m2_1312,m1[13],m2[12]);
and(m1m2_1313,m1[13],m2[13]);
and(m1m2_1314,m1[13],m2[14]);
and(m1m2_1315,m1[13],m2[15]);
and(m1m2_140,m1[14],m2[0]);
and(m1m2_141,m1[14],m2[1]);
and(m1m2_142,m1[14],m2[2]);
and(m1m2_143,m1[14],m2[3]);
and(m1m2_144,m1[14],m2[4]);
and(m1m2_145,m1[14],m2[5]);
and(m1m2_146,m1[14],m2[6]);
and(m1m2_147,m1[14],m2[7]);
and(m1m2_148,m1[14],m2[8]);
and(m1m2_149,m1[14],m2[9]);
and(m1m2_1410,m1[14],m2[10]);
and(m1m2_1411,m1[14],m2[11]);
and(m1m2_1412,m1[14],m2[12]);
and(m1m2_1413,m1[14],m2[13]);
and(m1m2_1414,m1[14],m2[14]);
and(m1m2_1415,m1[14],m2[15]);
and(m1m2_150,m1[15],m2[0]);
and(m1m2_151,m1[15],m2[1]);
and(m1m2_152,m1[15],m2[2]);
and(m1m2_153,m1[15],m2[3]);
and(m1m2_154,m1[15],m2[4]);
and(m1m2_155,m1[15],m2[5]);
and(m1m2_156,m1[15],m2[6]);
and(m1m2_157,m1[15],m2[7]);
and(m1m2_158,m1[15],m2[8]);
and(m1m2_159,m1[15],m2[9]);
and(m1m2_1510,m1[15],m2[10]);
and(m1m2_1511,m1[15],m2[11]);
and(m1m2_1512,m1[15],m2[12]);
and(m1m2_1513,m1[15],m2[13]);
and(m1m2_1514,m1[15],m2[14]);
and(m1m2_1515,m1[15],m2[15]);
buf(M[0],m1m2_00);
assign p0={1'b0,m1m2_150,m1m2_140,m1m2_130,m1m2_120,m1m2_110,m1m2_100,m1m2_90,m1m2_80,m1m2_70,m1m2_60,m1m2_50,m1m2_40,m1m2_30,m1m2_20,m1m2_10};
assign p1={m1m2_151,m1m2_141,m1m2_131,m1m2_121,m1m2_111,m1m2_101,m1m2_91,m1m2_81,m1m2_71,m1m2_61,m1m2_51,m1m2_41,m1m2_31,m1m2_21,m1m2_11,m1m2_01};
assign p2={m1m2_152,m1m2_142,m1m2_132,m1m2_122,m1m2_112,m1m2_102,m1m2_92,m1m2_82,m1m2_72,m1m2_62,m1m2_52,m1m2_42,m1m2_32,m1m2_22,m1m2_12,m1m2_02};
assign p3={m1m2_153,m1m2_143,m1m2_133,m1m2_123,m1m2_113,m1m2_103,m1m2_93,m1m2_83,m1m2_73,m1m2_63,m1m2_53,m1m2_43,m1m2_33,m1m2_23,m1m2_13,m1m2_03};
assign p4={m1m2_154,m1m2_144,m1m2_134,m1m2_124,m1m2_114,m1m2_104,m1m2_94,m1m2_84,m1m2_74,m1m2_64,m1m2_54,m1m2_44,m1m2_34,m1m2_24,m1m2_14,m1m2_04};
assign p5={m1m2_155,m1m2_145,m1m2_135,m1m2_125,m1m2_115,m1m2_105,m1m2_95,m1m2_85,m1m2_75,m1m2_65,m1m2_55,m1m2_45,m1m2_35,m1m2_25,m1m2_15,m1m2_05};
assign p6={m1m2_156,m1m2_146,m1m2_136,m1m2_126,m1m2_116,m1m2_106,m1m2_96,m1m2_86,m1m2_76,m1m2_66,m1m2_56,m1m2_46,m1m2_36,m1m2_26,m1m2_16,m1m2_06};
assign p7={m1m2_157,m1m2_147,m1m2_137,m1m2_127,m1m2_117,m1m2_107,m1m2_97,m1m2_87,m1m2_77,m1m2_67,m1m2_57,m1m2_47,m1m2_37,m1m2_27,m1m2_17,m1m2_07};
assign p8={m1m2_158,m1m2_148,m1m2_138,m1m2_128,m1m2_118,m1m2_108,m1m2_98,m1m2_88,m1m2_78,m1m2_68,m1m2_58,m1m2_48,m1m2_38,m1m2_28,m1m2_18,m1m2_08};
assign p9={m1m2_159,m1m2_149,m1m2_139,m1m2_129,m1m2_119,m1m2_109,m1m2_99,m1m2_89,m1m2_79,m1m2_69,m1m2_59,m1m2_49,m1m2_39,m1m2_29,m1m2_19,m1m2_09};
assign p10={m1m2_1510,m1m2_1410,m1m2_1310,m1m2_1210,m1m2_1110,m1m2_1010,m1m2_910,m1m2_810,m1m2_710,m1m2_610,m1m2_510,m1m2_410,m1m2_310,m1m2_210,m1m2_110,m1m2_010};
assign p11={m1m2_1511,m1m2_1411,m1m2_1311,m1m2_1211,m1m2_1111,m1m2_1011,m1m2_911,m1m2_811,m1m2_711,m1m2_611,m1m2_511,m1m2_411,m1m2_311,m1m2_211,m1m2_111,m1m2_011};
assign p12={m1m2_1512,m1m2_1412,m1m2_1312,m1m2_1212,m1m2_1112,m1m2_1012,m1m2_912,m1m2_812,m1m2_712,m1m2_612,m1m2_512,m1m2_412,m1m2_312,m1m2_212,m1m2_112,m1m2_012};
assign p13={m1m2_1513,m1m2_1413,m1m2_1313,m1m2_1213,m1m2_1113,m1m2_1013,m1m2_913,m1m2_813,m1m2_713,m1m2_613,m1m2_513,m1m2_413,m1m2_313,m1m2_213,m1m2_113,m1m2_013};
assign p14={m1m2_1514,m1m2_1414,m1m2_1314,m1m2_1214,m1m2_1114,m1m2_1014,m1m2_914,m1m2_814,m1m2_714,m1m2_614,m1m2_514,m1m2_414,m1m2_314,m1m2_214,m1m2_114,m1m2_014};
assign p15={m1m2_1515,m1m2_1415,m1m2_1315,m1m2_1215,m1m2_1115,m1m2_1015,m1m2_915,m1m2_815,m1m2_715,m1m2_615,m1m2_515,m1m2_415,m1m2_315,m1m2_215,m1m2_115,m1m2_015};
adder_16bit add0(p0,p1,1'b0,sum1,c1);
buf(M[1],sum1[0]);
adder_16bit add2({c1,sum1[15:1]},p2,1'b0,sum2,c2);
buf(M[2],sum2[0]);
adder_16bit add3({c2,sum2[15:1]},p3,1'b0,sum3,c3);
buf(M[3],sum3[0]);
adder_16bit add4({c3,sum3[15:1]},p4,1'b0,sum4,c4);
buf(M[4],sum4[0]);
adder_16bit add5({c4,sum4[15:1]},p5,1'b0,sum5,c5);
buf(M[5],sum5[0]);
adder_16bit add6({c5,sum5[15:1]},p6,1'b0,sum6,c6);
buf(M[6],sum6[0]);
adder_16bit add7({c6,sum6[15:1]},p7,1'b0,sum7,c7);
buf(M[7],sum7[0]);
adder_16bit add8({c7,sum7[15:1]},p8,1'b0,sum8,c8);
buf(M[8],sum8[0]);
adder_16bit add9({c8,sum8[15:1]},p9,1'b0,sum9,c9);
buf(M[9],sum9[0]);
adder_16bit add10({c9,sum9[15:1]},p10,1'b0,sum10,c10);
buf(M[10],sum10[0]);
adder_16bit add11({c10,sum10[15:1]},p11,1'b0,sum11,c11);
buf(M[11],sum11[0]);
adder_16bit add12({c11,sum11[15:1]},p12,1'b0,sum12,c12);
buf(M[12],sum12[0]);
adder_16bit add13({c12,sum12[15:1]},p13,1'b0,sum13,c13);
buf(M[13],sum13[0]);
adder_16bit add14({c13,sum13[15:1]},p14,1'b0,sum14,c14);
buf(M[14],sum14[0]);
adder_16bit add15({c14,sum14[15:1]},p15,1'b0,sum15,c15);
buf(M[15],sum15[0]);
assign out={sum15[0],M[14:0]};
endmodule